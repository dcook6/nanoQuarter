/*
* 	Derek Cook
* 	Minion CPU - NanoQuarter
*
*	Module:  Branch Adder TB
*	Inputs:  boff, PC_n, bne
*	Outputs: bse1
*
*/
module Branch_Adder_TB();

	reg[4:0] 	boff;
	reg[15:0]   	PC_n;
	reg         	bne;
	
	wire[15:0] 	bsel; 

	

	Branch_Adder test(.boff(boff), .PC_n(PC_n), .bne(bne), .bsel(bsel));


	initial begin
		
		#10 PC_n = 16'b0000000000000000;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000001;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000010;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000011;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000100;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000101;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000110;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000111;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001000;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001001;	bne = 0; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000000;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000001;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000010;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000011;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000100;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000101;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000110;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000111;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001000;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001001;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001010;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001100;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000001101;	bne = 1; boff = 4'b0000;
		#10 PC_n = 16'b0000000000000000;	bne = 1; boff = 4'b0001;
		#10 PC_n = 16'b0000000000000001;	bne = 1; boff = 4'b0010;
		#10 PC_n = 16'b0000000000000010;	bne = 1; boff = 4'b0011;
		#10 PC_n = 16'b0000000000000011;	bne = 1; boff = 4'b0100;
		#10 PC_n = 16'b0000000000000100;	bne = 1; boff = 4'b0101;
		#10 PC_n = 16'b0000000000000101;	bne = 1; boff = 4'b0110;
		#10 PC_n = 16'b0000000000000110;	bne = 1; boff = 4'b0111;
		#10 PC_n = 16'b0000000000000111;	bne = 1; boff = 4'b1000;
		#10 PC_n = 16'b0000000000001000;	bne = 1; boff = 4'b1001;
		#10 PC_n = 16'b0000000000001001;	bne = 1; boff = 4'b1010;
		#10 PC_n = 16'b0000000000001010;	bne = 1; boff = 4'b1011;
		#10 PC_n = 16'b0000000000001100;	bne = 1; boff = 4'b1100;
		#10 PC_n = 16'b0000000000001101;	bne = 1; boff = 4'b1111;
		#10 PC_n = 16'b0000000000000000;	bne = 0; boff = 4'b0001;
		#10 PC_n = 16'b0000000000000001;	bne = 0; boff = 4'b0010;
		#10 PC_n = 16'b0000000000000010;	bne = 0; boff = 4'b0011;
		#10 PC_n = 16'b0000000000000011;	bne = 0; boff = 4'b0100;
		#10 PC_n = 16'b0000000000000100;	bne = 0; boff = 4'b0101;
		#10 PC_n = 16'b0000000000000101;	bne = 0; boff = 4'b0110;
		#10 PC_n = 16'b0000000000000110;	bne = 0; boff = 4'b0111;
		#10 PC_n = 16'b0000000000000111;	bne = 0; boff = 4'b1000;
		#10 PC_n = 16'b0000000000001000;	bne = 0; boff = 4'b1001;
		#10 PC_n = 16'b0000000000001001;	bne = 0; boff = 4'b1010;
		#10 PC_n = 16'b0000000000001010;	bne = 0; boff = 4'b1011;
		#10 PC_n = 16'b0000000000001100;	bne = 0; boff = 4'b1100;
		#10 PC_n = 16'b0000000000001101;	bne = 0; boff = 4'b1111;		
		$finish;

	end
endmodul
